library ieee;
use ieee.std_logic_1164.all;

--constants, components, 
package test_pkg is
	--constant declaration
	constant NAME : integer := 720;
end package;


