library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.math_pkg.all;

use work.test_pkg.all;

-- TODO: add entity (generic: constants, ports: inputs/outputs)
entity design_name is
end entity;

-- TODO: add implementation of design
architecture beh of design_name is 
-- TODO: add signals, declare-components
begin 
	-- TODO: add design (process, concurrent-statements, init-components)
end architecture;