library ieee;
use ieee.std_logic_1164.all;

package test_pkg is
	constant NAME : integer := 720;
end package;


