library ieee;
use ieee.std_logic_1164.all;

package helper_pkg is 
	constant SCREEN_WIDTH_TEST : natural := 300;

	--define components 
end package;