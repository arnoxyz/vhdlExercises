library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.math_pkg.all;
use work.test_pkg.all;


--simple_timer
entity simple_timer is

end entity;


--FSM Template 
--simple timer

architecture arch of simple_timer is 
begin 
end architecture;
