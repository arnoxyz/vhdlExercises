library ieee;
use ieee.std_logic_1164.all;

--define some constants that can be used in the design
package test_pkg is
	--constant declaration
	constant SCREEN_WIDTH : integer := 720;
	constant SCREEN_HEIGHT : integer := 480;
end package;


